module test;
    initial $display("%0b", 1'b1 | 4'b1010);
endmodule