module test;
    initial $display("%0b", 4'b1010 & 4'b1000);
endmodule