module signed_cmp_;
endmodule