module integer_issue_golden #() (

);
    // state elements
    