module dff_we();

endmodule