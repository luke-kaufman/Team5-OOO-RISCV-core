module load_store_execute #(

) (
    input wire clk,
    input wire rst_aL,

);
    
endmodule