// IMPL STATUS: MISSING
// TEST STATUS: MISSING
module onehot_mux4 (
    input wire [3:0] sel,
    input wire [3:0] din,
    output wire dout
);
endmodule