module memory(
    input [31:0] address_bus,
    inout [31:0] data_bus,
    input read,
    input write
    );

endmodule