module test;
    $display("%0b", 4'b1010 & 1'b1);
endmodule