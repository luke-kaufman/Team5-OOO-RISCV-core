module top(
);



endmodule