module ifu(
    output wire [:] inst_o;
    
);

endmodule