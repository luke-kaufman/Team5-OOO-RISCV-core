module predicted_NPC # (

) (

);
endmodule