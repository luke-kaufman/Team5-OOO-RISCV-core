module RAT #() (

);
    Regfile #() arf_rob (

    );

    Regfile #() 

endmodule