`include "misc/global_defs.svh"
`include "top/top.sv"

module dispatch_tb #(
    parameter addr_t HIGHEST_PC = 32'h1018c,
    localparam main_mem_block_addr_t HIGHEST_INSTR_BLOCK_ADDR = HIGHEST_PC >> `MAIN_MEM_BLOCK_OFFSET_WIDTH
);
    bit clk = 0;
    bit init = 0;
    addr_t init_pc = 32'h1018c;
    addr_t init_sp = init_pc - 4;
    main_mem_block_addr_t block_addr;
    main_mem_block_offset_t block_offset;
    // block_data_t init_main_mem_state[`MAIN_MEM_N_BLOCKS];
    block_data_t init_main_mem_state[HIGHEST_INSTR_BLOCK_ADDR:0];

    initial forever #5 clk = ~clk;

    initial begin
        // for (int i = 0; i < `MAIN_MEM_N_BLOCKS; i++) begin // TODO: double-check if this is correct
        //     init_main_mem_state[i] = '0;
        // end
        {block_addr, block_offset} = 32'h1018c; // 0001 0000 0001 1000 1100
        if (8*block_offset + `INSTR_WIDTH <= `BLOCK_DATA_WIDTH) begin
            // init_main_mem_state[block_addr][8*block_offset+:`INSTR_WIDTH] = 32'hfe010113;
            init_main_mem_state[HIGHEST_INSTR_BLOCK_ADDR][8*block_offset+:`INSTR_WIDTH] = 32'hfe010113;
        end
        // else begin
        //     automatic logic [`BLOCK_DATA_WIDTH-block_offset-1:0] instr_part1;
        //     automatic logic [`INSTR_WIDTH-$bits(instr_part1)-1:0] instr_part2;
        //     {instr_part1, instr_part2} = 32'hfe010113;
        //     init_main_mem_state[block_addr][`BLOCK_DATA_WIDTH-1:block_offset] = instr_part1;
        //     init_main_mem_state[block_addr+1][$bits(instr_part2)-1:0] = instr_part2;
        // end
    end


    wire [`ARF_N_ENTRIES-1:0] [`REG_DATA_WIDTH-1:0] ARF_OUT;

    top #(
        .HIGHEST_PC(HIGHEST_PC)
    ) _top (
        .clk(clk),
        .rst_aL(),
        .init(init),
        .init_pc(init_pc),
        .init_sp(init_sp),
        .init_main_mem_state(init_main_mem_state),
        .ARF_OUT(ARF_OUT)
    );

    initial begin
        // $display("%0t way1_data: %b", $time, _top._core._ifu.icache.data_array_dout.way1_data);
        #101 $display("%0t way1_data: %b", $time, _top._core._ifu.icache.data_array_dout.way1_data);

        $display("%0t sel_data_behind[0]: %b", $time, _top._core.integer_issue_dut.iiq.sel_data_behind[0]);
        $display("%0t sel_enq_data[0]: %b", $time, _top._core.integer_issue_dut.iiq.sel_enq_data[0]);
        $display("%0t sel_wr_data[0]: %b", $time, _top._core.integer_issue_dut.iiq.sel_wr_data[0]);
        $display("%0t sel_wr_data_behind[0]: %b", $time, _top._core.integer_issue_dut.iiq.sel_wr_data_behind[0]);
    end

    initial begin
        // $monitor("%b", ARF_OUT);
        $monitor("%0t PC_mux_out: %b", $time, _top._core._ifu.PC_mux_out);
        $monitor("%0t ififo: %h", $time, _top._core._ifu.instruction_FIFO);

        // $monitor("%p", _top._main_mem.mem);
        // $monitor("%b", _top._mem_ctrl.icache_req_valid);
        // $monitor("%b", _top._mem_ctrl.icache_req_block_addr);
        // $monitor("%b", _top._mem_ctrl.icache_req_ready);
        // $monitor("%t, %p", $time, _top._main_mem.req_pipeline);

        #1;
        init = 1;
        #1;
        init = 0;
        #1;
        @(negedge clk);
        @(negedge clk);
        repeat (10)
            @(negedge clk);
        $finish;
    end
endmodule
