// IMPL STATUS: MISSING
// TEST STATUS: MISSING
module mux2 #(
    parameter WIDTH = 1
) (
    input wire sel,
    input wire [WIDTH-1:0] in0,
    input wire [WIDTH-1:0] in1,
    output wire [WIDTH-1:0] out
);

endmodule