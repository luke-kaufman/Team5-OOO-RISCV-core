module load_store_issue #(

) (

);
    shift_queue lsq (
        // .clk(clk),
        // .rst_aL(rst_aL),
        // .enq_ready(),
        // .enq_valid(),
        // .enq_data(),
        // .deq_ready(),
        // .deq_valid(),
        // .deq_data()
    );
endmodule