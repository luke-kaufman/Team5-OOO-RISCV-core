module icache_data_bank (
    input wire clk,
    input wire rst
    
);
    
endmodule