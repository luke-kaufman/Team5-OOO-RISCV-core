module icache_tag_bank #(
    parameter WORD_SIZE = 32,
    parameter N_WORDS = 64
) (
    input wire clk,
    input wire rst,
    input wire en,
    output wire [WORD_SIZE-1:0] dout
);
    
endmodule