`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/28/2024 06:03:20 PM
// Design Name: 
// Module Name: ADDER_EN_32in
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ADDER_EN_32in(
    input[31:0] in1, in2,
    output[31:0] data_out
    );
    assign data_out = in1 + in2;
endmodule
