`ifndef SHIFT_QUEUE_V
`define SHIFT_QUEUE_V

`include "misc/reg_.v"
`include "misc/up_down_counter.v"
`include "misc/cmp/unsigned_cmp_.v"
`include "misc/onehot_mux/onehot_mux_.v"
`include "misc/dec/dec_.v"
`include "misc/and/and_.v"
`include "misc/or/or_.v"
`include "misc/extend_first1.v"

// IMPL STATUS: COMPLETE
// TEST STATUS: MISSING
module shift_queue #(
    parameter N_ENTRIES = `IIQ_N_ENTRIES,
    parameter ENTRY_WIDTH = `IIQ_ENTRY_WIDTH,
    localparam PTR_WIDTH = $clog2(N_ENTRIES),
    localparam CTR_WIDTH = PTR_WIDTH + 1
) (
    input wire clk,
    input wire rst_aL,

    // enqueue interface: ready & valid
    output wire enq_ready,
    input wire enq_valid,
    input wire [ENTRY_WIDTH-1:0] enq_data,

    // dequeue interface: select then valid
    input wire deq_ready,
    input wire [N_ENTRIES-1:0] deq_sel_onehot, // can be either one-hot or all 0s
    output wire deq_valid,
    output wire [ENTRY_WIDTH-1:0] deq_data,

    input wire [N_ENTRIES-1:0] wr_en,
    input wire [N_ENTRIES-1:0] [ENTRY_WIDTH-1:0] wr_data,

    output wire [N_ENTRIES-1:0] [ENTRY_WIDTH-1:0] entry_douts,
    output wire [CTR_WIDTH-1:0] enq_ctr_dout,

    input wire flush,

    // for testing
    input wire init,
    input wire [N_ENTRIES-1:0] [ENTRY_WIDTH-1:0] init_entry_reg_state,
    input wire [CTR_WIDTH-1:0] init_enq_up_down_counter_state,
    output wire [N_ENTRIES-1:0] [ENTRY_WIDTH-1:0] current_entry_reg_state,
    output wire [CTR_WIDTH-1:0] current_enq_up_down_counter_state
);
    // internal signal
    wire [CTR_WIDTH-1:0] enq_ctr; // one bit wider than the pointer width to allow for the full condition (we can still enqueue to the queue when it is full if there will be a dequeue in the same cycle)
    wire [PTR_WIDTH-1:0] enq_ptr = enq_ctr[PTR_WIDTH-1:0]; // the enqueue pointer is the lower bits of the enqueue counter
    wire queue_full = enq_ctr[PTR_WIDTH]; // the queue is full if the MSB of the enqueue counter is true
    wire enq;
    and_ #(.N_INS(2)) enq_and (
        .a({enq_ready, enq_valid}),
        .y(enq)
    );
    wire deq;
    and_ #(.N_INS(2)) deq_and (
        .a({deq_ready, deq_valid}),
        .y(deq)
    );
    // extend the dequeue select signal to generate the precursor write enable signals generated by the dequeue interface
    wire [N_ENTRIES-1:0] shift_we_pre;
    extend_first1 #(.WIDTH(N_ENTRIES)) shift_we_pre_extf1 (
        .a(deq_sel_onehot),
        .y(shift_we_pre)
    );
    // gate the shift_we_pre signal with the dequeue signal so that the shift_we signal is only true when the dequeue signal is true
    wire [N_ENTRIES-1:0] shift_we;
    for (genvar i = 0; i < N_ENTRIES; i++) begin
        and_ #(.N_INS(2)) shift_we_and (
            .a({shift_we_pre[i], deq}),
            .y(shift_we[i])
        );
    end
    wire [N_ENTRIES:0] enq_we_ext_pre;
    wire [2**CTR_WIDTH-1:0] enq_ctr_decoder_out;
    // decode the enqueue pointer (lower bits of the enqueue counter) to generate the precursor extended write enable signals generated by the enqueue interface
    dec_ #(.IN_WIDTH(CTR_WIDTH)) enq_ctr_decoder (
        .in(enq_ctr),
        .out(enq_ctr_decoder_out)
    );
    assign enq_we_ext_pre = enq_ctr_decoder_out[N_ENTRIES:0]; // the (one-hot) enqueue write enable signal is the lower bits of the decoder output

    // gate the enq_we_ext_pre signal with the enqueue signal so that the enq_we_ext signal is only true when the enqueue signal is true
    wire [N_ENTRIES:0] enq_we_ext;
    for (genvar i = 0; i <= N_ENTRIES; i++) begin
        and_ #(.N_INS(2)) enq_we_and (
            .a({enq_we_ext_pre[i], enq}),
            .y(enq_we_ext[i])
        );
    end

    wire [N_ENTRIES:0] wr_en_ext = {1'b0, wr_en}; // write enable extended (last element is false because the outside of the queue can't be written to)

    // the events dequeue and shift are if and only if conditions (i.e. dequeue is true iff shift is true)
    // the concrete examples of enqueue, dequeue, and write signals in this formulation, for the case of integer issue queue:
    // - enqueue = dispatch
    // - dequeue (= shift) = issue
    // - write = wakeup
    // write and shift case:
    // - the write data is shifted as well (register i-1 gets the write data, register i doesn't) (NOTE: writes to register 0 don't shift)
    // enqueue and shift case:
    // - the enqueued entry is shifted as well (register i-1 gets the enqueued entry, register i doesn't) (NOTE: enqueues to register 0 don't shift)
    // so, the (one-hot) din_mux of register i chooses between:
    // - enq_data (if enq is true AND (shift is true AND enq_we_ext[i+1] is true OR shift is false AND enq_ptr[i] is true)) (NOTE: enq_we_ext[i+1] exists even for i = N_ENTRIES-1)
    // - wr_data (if wr_en[i] is true AND shift is false OR wr_en[i+1] is true AND shift is true) (NOTE: wr_en[i+1] is 1'b0 instead for i = N_ENTRIES-1 (there won't be a write to outside of the queue))
    // - entry_douts[i+1] (if shift is true) (NOTE: entry_douts[i+1] is {ENTRY_WIDTH{1'b0}} instead if i = N_ENTRIES-1)
    // shift_we[i] | enq_we_ext[i+1] | wr_en[i+1] | enq_we_ext[i] | wr_en[i] | din[i]
    // 0           | x               | x          | 0             | 0        | entry_douts[i]
    // 0           | x               | x          | 0             | 1        | wr_data[i]
    // 0           | x               | x          | 1             | 0        | enq_data
    // 0           | x               | x          | 1             | 1        | error (we cannot write to empty entries)
    // 1           | 0               | 0          | x             | x        | entry_douts[i+1] (or {ENTRY_WIDTH{1'b0}} if i = N_ENTRIES-1)
    // 1           | 0               | 1          | x             | x        | wr_data[i+1] (or 1'b0 for i = N_ENTRIES-1)
    // 1           | 1               | 0          | x             | x        | enq_data
    // 1           | 1               | 1          | x             | x        | error (we cannot write to empty entries)
    // the select signals are generated by the following inputs:
    // - shift_we[i]
    // - wr_en_ext[i]
    // - enq_we_ext[i]
    // - wr_en_ext[i+1] (is 0 for i = N_ENTRIES-1)
    // - enq_we_ext[i+1] (exists even for i = N_ENTRIES-1)
    // so, the (one-hot) din_mux of register i chooses between:
    // - 0: entry_douts[i+1] (if shift_we[i] is true AND enq_we_ext[i+1] is false AND wr_en_ext[i+1] is false) (is all 0s if i = N_ENTRIES-1)
    // - 1: enq_data (if shift_we[i] is false and enq_we_ext[i] is true OR shift_we[i] is true and enq_we_ext[i+1] is true)
    // - 2: wr_data[i] (if shift_we[i] is false and wr_en_ext[i] is true)
    // - 3: wr_data[i+1] (if shift_we[i] is true and wr_en_ext[i+1] is true)
    // - default: if all the above conditions are false, register i should hold the same value as before
    // since we of register i is false anyway, the output of the mux is don't care (physically all 0s because of the one-hot mux implementation)
    // sel[0] = shift_we[i] & ~enq_we_ext[i+1] & ~wr_en_ext[i+1]
    // sel[1] = ~shift_we[i] & enq_we_ext[i] | shift_we[i] & enq_we_ext[i+1]
    // sel[2] = ~shift_we[i] & wr_en_ext[i]
    // sel[3] = shift_we[i] & wr_en_ext[i+1]
    wire [N_ENTRIES-1:0] shift_we_not;
    wire [N_ENTRIES:0] enq_we_ext_not;
    wire [N_ENTRIES:0] wr_en_ext_not;
    for (genvar i = 0; i < N_ENTRIES; i++) begin
        INV_X1 shift_we_inv (
            .A(shift_we[i]),
            .ZN(shift_we_not[i])
        );
        INV_X1 enq_we_ext_inv (
            .A(enq_we_ext[i]),
            .ZN(enq_we_ext_not[i])
        );
        INV_X1 wr_en_ext_inv (
            .A(wr_en_ext[i]),
            .ZN(wr_en_ext_not[i])
        );
    end
    INV_X1 enq_we_ext_last_inv (
        .A(enq_we_ext[N_ENTRIES]),
        .ZN(enq_we_ext_not[N_ENTRIES])
    );
    INV_X1 wr_en_ext_last_inv (
        .A(wr_en_ext[N_ENTRIES]),
        .ZN(wr_en_ext_not[N_ENTRIES])
    );

    //
    wire [N_ENTRIES-1:0] sel_data_behind; // sel[0]: entry_douts[i+1]
    for (genvar i = 0; i < N_ENTRIES; i++) begin
        and_ #(.N_INS(3)) sel_data_behind_and (
            .a({shift_we[i], enq_we_ext_not[i+1], wr_en_ext_not[i+1]}),
            .y(sel_data_behind[i])
        );
    end
    //

    //
    wire [N_ENTRIES-1:0] sel_enq_data_pre_from_this; // sel[1] -- ~shift_we[i] & enq_we_ext[i]
    wire [N_ENTRIES-1:0] sel_enq_data_pre_from_behind; // sel[1] -- shift_we[i] & enq_we_ext[i+1]
    wire [N_ENTRIES-1:0] sel_enq_data; // sel[1]: enq_data
    for (genvar i = 0; i < N_ENTRIES; i++) begin
        and_ #(.N_INS(2)) sel_enq_data_pre_from_this_and (
            .a({enq_we_ext[i], shift_we_not[i]}),
            .y(sel_enq_data_pre_from_this[i])
        );
        and_ #(.N_INS(2)) sel_enq_data_pre_from_behind_and (
            .a({enq_we_ext[i+1], shift_we[i]}),
            .y(sel_enq_data_pre_from_behind[i])
        );
        or_ #(.N_INS(2)) sel_enq_data_or (
            .a({sel_enq_data_pre_from_this[i], sel_enq_data_pre_from_behind[i]}),
            .y(sel_enq_data[i])
        );
    end
    //

    //
    wire [N_ENTRIES-1:0] sel_wr_data; // sel[2]: wr_data[i]
    for (genvar i = 0; i < N_ENTRIES; i++) begin
        and_ #(.N_INS(2)) sel_wr_data_and (
            .a({wr_en_ext[i], shift_we_not[i]}),
            .y(sel_wr_data[i])
        );
    end
    //

    //
    wire [N_ENTRIES-1:0] sel_wr_data_behind; // sel[3]: wr_data[i+1]
    for (genvar i = 0; i < N_ENTRIES; i++) begin
        and_ #(.N_INS(2)) sel_wr_data_behind_and (
            .a({wr_en_ext[i+1], shift_we[i]}),
            .y(sel_wr_data_behind[i])
        );
    end
    //

    // if wr_en_ext is true for empty entries (entries i where i >= enq_ptr), then throw an error TODO
    // assert(!|wr_en[N_ENTRIES-1:enq_ptr]|) else $fatal(0, "shift_queue: wr_en_ext is true for empty entries");

    // if all select signals are zero, the output is don't care (physically 0); the entry_we for the register is false anyway
    wire [N_ENTRIES-1:0] [ENTRY_WIDTH-1:0] entry_din;
    for (genvar i = 0; i < N_ENTRIES-1; i++) begin
        onehot_mux_ #(.WIDTH(ENTRY_WIDTH), .N_INS(4)) entry_din_mux (
            .clk(clk),
            .ins({entry_douts[i+1], enq_data, wr_data[i], wr_data[i+1]}),
            .sel({sel_data_behind[i], sel_enq_data[i], sel_wr_data[i], sel_wr_data_behind[i]}),
            .out(entry_din[i])
        );
    end
    onehot_mux_ #(.WIDTH(ENTRY_WIDTH), .N_INS(4)) entry_din_last_mux (
        // if sel_data_behind[N_ENTRIES-1] is true, then shift in fresh all 0s
        // sel_wr_data_behind[N_ENTRIES-1] is always false anyway
        .clk(clk),
        .ins({{ENTRY_WIDTH{1'b0}}, enq_data, wr_data[N_ENTRIES-1], {ENTRY_WIDTH{1'b0}}}),
        .sel({sel_data_behind[N_ENTRIES-1], sel_enq_data[N_ENTRIES-1], sel_wr_data[N_ENTRIES-1], sel_wr_data_behind[N_ENTRIES-1]}),
        .out(entry_din[N_ENTRIES-1])
    );

    // combine the select signals to generate the write enable signals for each entry
    wire [N_ENTRIES-1:0] entry_we;
    for (genvar i = 0; i < N_ENTRIES; i++) begin
        or_ #(.N_INS(4)) entry_we_or (
            .a({sel_data_behind[i], sel_enq_data[i], sel_wr_data[i], sel_wr_data_behind[i]}),
            .y(entry_we[i])
        );
    end

    // TODO: redundant with the implementation of up_down_counter (it already handles the case inc = 1, dec = 1)
    wire enq_ctr_inc;
    wire enq_ctr_dec;
    wire enq_not;
    wire deq_not;
    INV_X1 enq_inv (
        .A(enq),
        .ZN(enq_not)
    );
    INV_X1 deq_inv (
        .A(deq),
        .ZN(deq_not)
    );
    and_ #(.N_INS(2)) enq_ctr_inc_and (
        .a({enq, deq_not}),
        .y(enq_ctr_inc)
    );
    and_ #(.N_INS(2)) enq_ctr_dec_and (
        .a({enq_not, deq}),
        .y(enq_ctr_dec)
    );

    // output drivers
    // if the queue is not full OR there will be a dequeue, then enq_ready is true
    // WARNING: with this implementation, now the enqueue interface depends on the dequeue interface
    // TODO: check this for feasibility
    wire queue_not_full;
    INV_X1 inv (
        .A(queue_full),
        .ZN(queue_not_full)
    );
    or_ #(.N_INS(2)) enq_ready_or (
        .a({queue_not_full, deq}),
        .y(enq_ready)
    );

    // if any entry is selected for dequeue, then deq_valid is true
    or_ #(.N_INS(N_ENTRIES)) deq_valid_or (
        .a(deq_sel_onehot),
        .y(deq_valid)
    );
    // select the entry to be dequeued (outputs {ENTRY_WIDTH{1'b0}} when no entry is selected)
    onehot_mux_ #(.WIDTH(ENTRY_WIDTH), .N_INS(N_ENTRIES)) deq_data_mux (
        .clk(clk),
        .sel(deq_sel_onehot),
        .ins(entry_douts),
        .out(deq_data)
    );
    // entry_douts is already driven in each entry_reg instantiation

    // state elements
    up_down_counter #(.WIDTH(CTR_WIDTH)) enq_up_down_counter ( // NOTE: STATEFUL
        .clk(clk),
        .rst_aL(rst_aL),
        .inc(enq_ctr_inc),
        .dec(enq_ctr_dec),
        .count(enq_ctr),
        .flush(flush),
        .init(init),
        .init_state(init_enq_up_down_counter_state)
    );
    assign enq_ctr_dout = enq_ctr;
    for (genvar i = 0; i < N_ENTRIES; i++) begin : queue
        reg_ #(.WIDTH(ENTRY_WIDTH)) entry_reg ( // NOTE: STATEFUL
            .flush(flush),
            .clk(clk),
            .rst_aL(rst_aL),
            .we(entry_we[i]),
            .din(entry_din[i]),
            .dout(entry_douts[i]),

            .init(init),
            .init_state(init_entry_reg_state[i])
        );
    end

    assign current_entry_reg_state = entry_douts;
    assign current_enq_up_down_counter_state = enq_ctr;

    // assertions
    function void enq_ctr_max_value(edge_t _edge);
        if (enq_ctr > N_ENTRIES) begin
            $error(
                "%0t Assertion failed: enq_ctr is larger than max value after %0s.\n\
                enq_ctr = %0d, max value = %0d\n",
                $time, _edge == NEGEDGE ? "setting init_state and driving inputs" : "state transition",
                enq_ctr, N_ENTRIES
            );
            $display("%0t enq_valid: %b, enq_ready: %b, deq_ready: %b, deq_sel_onehot: %b, deq_valid: %b",
                    $time, enq_valid, enq_ready, deq_ready, deq_sel_onehot, deq_valid);
        end
    endfunction

    always @(negedge clk) begin #1
        enq_ctr_max_value(NEGEDGE);
    end
    always @(posedge clk) begin #1
        enq_ctr_max_value(POSEDGE);
    end
endmodule

`endif
