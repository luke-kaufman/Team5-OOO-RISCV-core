module core(
    input [31:0] address_bus,
    inout [31:0] data_bus,
    output memory_read,
    output memory_write
);

    

endmodule