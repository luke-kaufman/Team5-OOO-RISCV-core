// IMPL STATUS: MISSING
// TEST STATUS: MISSING
module ff1 (

);
endmodule