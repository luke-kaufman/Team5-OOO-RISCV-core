module load_store_issue #(

) (

);
    shift_queue lsq (
        // .clk(clk),
        // .rst_aL(rst_aL),
        // .ready_enq(),
        // .valid_enq(),
        // .data_enq(),
        // .ready_deq(),
        // .valid_deq(),
        // .data_deq()
    );
endmodule