module instruction_FIFO # (

) (

);

endmodule